module mul4 (s, a, b);
output [8:0] s;
input  [3:0] a, b;
assign s = a * b;
endmodule
